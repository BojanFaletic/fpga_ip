library ieee;
use ieee.std_logic_1164.all;

package image_generator_pkg is
  constant C_LINE_WIDTH : integer := 230;
  constant C_LINE_HEIGHT : integer := 355;
  constant C_IS_GRAY : boolean := False;
  constant C_FILENAME : string := "cat.coe";
end package;

package body image_generator_pkg is
end package body;